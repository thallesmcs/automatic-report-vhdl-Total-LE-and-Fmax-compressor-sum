library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity FF_D8 is
    port (
        clk   : in  std_logic;
        rst_n : in  std_logic;  -- reset assíncrono ativo baixo
        d     : in  std_logic_vector(7 downto 0);
        q     : out std_logic_vector(7 downto 0)
    );
end entity;

architecture rtl of FF_D8 is
begin
    process (clk, rst_n)
    begin
        if rst_n = '0' then          -- reset assíncrono ativo baixo
            q <= (others => '0');
        elsif rising_edge(clk) then
            q <= d;
        end if;
    end process;
end architecture;
